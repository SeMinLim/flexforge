import FIFO::*;
import FIFOF::*;
import Clocks::*;
import Vector::*;

import Serializer::*;

import BRAM::*;
import BRAMFIFO::*;

import PcieCtrl::*;

import DRAMController::*;
import DRAMArbiterRemote::*;

import Kmean::*;

Integer numData = 1024;
Integer totalByte = 2*1024*4;
Integer totalWords = 2*64;
Integer bramFifoSize = 1024;

typedef 1024 NumData;
typedef 4 PeWaysLog;
typedef TExp#(PeWaysLog) PeWays;


interface HwMainIfc;
endinterface
module mkHwMain#(PcieUserIfc pcie, DRAMUserIfc dram) (HwMainIfc);

	Clock curClk <- exposeCurrentClock;
	Reset curRst <- exposeCurrentReset;

	Clock pcieclk = pcie.user_clk;
	Reset pcierst = pcie.user_rst;

	// Cycle Counter
	FIFOF#(Bit#(32)) cycleQ <- mkFIFOF;
	Reg#(Bit#(32)) cycleCount <- mkReg(0);
	Reg#(Bit#(32)) cycleStart <- mkReg(0);
	Reg#(Bit#(32)) cycleEnd <- mkReg(0);
	rule incCycleCount;
		cycleCount <= cycleCount + 1;
	endrule

	// Serializer
	DeSerializerIfc#(32, 16) deserializer32b <- mkDeSerializer;
	SerializerIfc#(512, 8) serializer64b <- mkSerializer;

	// DRAM Arbiter
	DRAMArbiterRemoteIfc#(2) dramArbiter <- mkDRAMArbiterRemote(dram);
	
	// K-mean App
	KmeanIfc kmean <- mkKmean;
	//--------------------------------------------------------------------------------------
	// Pcie Read and Write
	//--------------------------------------------------------------------------------------
	SyncFIFOIfc#(Tuple2#(IOReadReq, Bit#(32))) pcieRespQ <- mkSyncFIFOFromCC(1024, pcieclk);
	SyncFIFOIfc#(IOReadReq) pcieReadReqQ <- mkSyncFIFOToCC(1024, pcieclk, pcierst);
	SyncFIFOIfc#(IOWrite) pcieWriteQ <- mkSyncFIFOToCC(1024, pcieclk, pcierst);
	rule getReadReq;
		let r <- pcie.dataReq;
		pcieReadReqQ.enq(r);
	endrule
	rule returnReadResp;
		let r_ = pcieRespQ.first;
		pcieRespQ.deq;

		pcie.dataSend(tpl_1(r_), tpl_2(r_));
	endrule
	rule getWriteReq;
		let w <- pcie.dataReceive;
		pcieWriteQ.enq(w);
	endrule
	//--------------------------------------------------------------------------------------------
	// Get Commands from Host via PCIe
	//--------------------------------------------------------------------------------------------
	FIFOF#(Bit#(32)) statusCheckerQ <- mkFIFOF;
	// Initial Setting
	Reg#(Bool) stage1 <- mkReg(False);
	// DRAM Reader
	Reg#(Bool) stage2 <- mkReg(False);
	// Data Serializer
	Reg#(Bool) stage3 <- mkReg(False);
	Reg#(Bool) enqClusterHeadQ <- mkReg(True);
	// Data Relayer
	Reg#(Bool) stage4 <- mkReg(False);
	// Data Receiver
	Reg#(Bool) stage5 <- mkReg(False);
	rule getCmd;
		pcieWriteQ.deq;
		let w = pcieWriteQ.first;

		let d = w.data;
		let a = w.addr;
		let off = (a >> 2);

		if ( off == 0 ) begin
			stage1 <= True;
			$write("\033[1;33mCycle %1d -> \033[1;33m[HwMain]: \033[0m: Initial setting start!\n", cycleCount);
		end else if ( off == 1 ) begin
			deserializer32b.put(d);
		end else if ( off == 2 ) begin
			stage2 <= True;
			stage3 <= True;
			stage4 <= True;
			stage5 <= True;
			$write("\033[1;33mCycle %1d -> \033[1;33m[HwMain]: \033[0m: System start!\n", cycleCount);
		end
	endrule
	//--------------------------------------------------------------------------------------------
	// Usage of the entire memory
	//  For Mode 1
	//  0 ~ 8,191
	//--------------------------------------------------------------------------------------------
	// Stage 1 (Initial Setting)
	//
	// This stage writes the data take from the host through PCIe to DRAM
	//--------------------------------------------------------------------------------------------
	Reg#(Bit#(32)) stage1Cnt <- mkReg(0); // Good!!!
	rule dramWriterInit( stage1 );
		if ( stage1Cnt != 0 ) begin
			let payload <- deserializer32b.get;
			dramArbiter.access[0].users[0].write(payload);
			if ( stage1Cnt == fromInteger(totalWords) ) begin
				stage1Cnt <= 0;
				stage1 <= False;

				//statusCheckerQ.enq(1); // Check dram writer initial set done
				$write("\033[1;33mCycle %1d -> \033[1;33m[HwMain]: \033[0m: Initial setting \033[1;32mdone!\n", cycleCount);
			end else begin
				stage1Cnt <= stage1Cnt + 1;
			end
		end else begin
			dramArbiter.access[0].users[0].cmd(0, fromInteger(totalWords), True);
			stage1Cnt <= stage1Cnt + 1;
		end
	endrule
	//--------------------------------------------------------------------------------------------
	// Stage 2 (DRAM Reader)
	//
	// This stage read the data from DRAM
	//--------------------------------------------------------------------------------------------
	Reg#(Bit#(16)) stage2Cnt <- mkReg(0); // Good!!!
	rule dramReader( stage2 );
		if ( stage2Cnt != 0 ) begin
			let payload <- dramArbiter.access[0].users[0].read;
			serializer64b.put(payload);
				
			if ( stage2Cnt == 128 ) begin
				stage2Cnt <= 0;
				$write("\033[1;33mCycle %1d -> \033[1;33m[HwMain]: \033[0m: Read 1024 x and y data \033[1;32mdone!\n", cycleCount);
				stage2 <= False;
			end else begin
				stage2Cnt <= stage2Cnt + 1;
			end
		end else begin
			dramArbiter.access[0].users[0].cmd(0, 128, False); // 2*1024*4 = 128*64
			stage2Cnt <= stage2Cnt + 1;
			$write("\033[1;33mCycle %1d -> \033[1;33m[HwMain]: \033[0m: Read 1024 x and y data \033[1;32mstart!\n", cycleCount);
		end
	endrule
	//-------------------------------------------------------------------------------------------------
	// Stage 3 (Data Serializer)
	//
	// This state splits the 512-bit payload to 32-bit data
	//-------------------------------------------------------------------------------------------------
	FIFO#(Vector#(2, Bit#(32))) originDataQ <- mkSizedBRAMFIFO(1024);
	FIFO#(Vector#(2, Bit#(32))) clusterHeadQ <- mkSizedBRAMFIFO(16);
	Reg#(Bit#(16)) stage3Cnt <- mkReg(0);
	Reg#(Bit#(16)) testCnt <- mkReg(0);
	rule dataSerializer( stage3 );
		Vector#(2, Bit#(32)) v = replicate(0);
		let d <- serializer64b.get;
		v[0] = d[31:0]; // x
		v[1] = d[63:32]; // y
		
		originDataQ.enq(v);
		
		if ( enqClusterHeadQ ) begin
			if ( stage3Cnt + 1 == fromInteger(valueOf(PeWays)) ) begin
				stage3Cnt <= 0;
				enqClusterHeadQ <= False;
			end else begin
				stage3Cnt <= stage3Cnt + 1;
			end
			clusterHeadQ.enq(v);
		end
	endrule
	//--------------------------------------------------------------------------------------------
	// Stage 4 (K-mean, Data Relayer)
	//
	// This stage relays the data to K-mean app
	//--------------------------------------------------------------------------------------------
	Reg#(Bit#(16)) stage4Cnt_1 <- mkReg(0);
	rule dataRelayer( stage4 );
		originDataQ.deq;
		let v = originDataQ.first;

		kmean.dataIn(v);

		if ( stage4Cnt_1 + 1 == fromInteger(bramFifoSize) ) begin
			stage4Cnt_1 <= 0;
			$write("\033[1;33mCycle %1d -> \033[1;33m[HwMain]: \033[0m: Relay 1024 x and y data \033[1;32mdone!\n", cycleCount);
		end else begin
			stage4Cnt_1 <= stage4Cnt_1 + 1;
		end
	endrule

	Reg#(Bit#(16)) stage4Cnt_2 <- mkReg(0);
	rule dataRelayer_ClusterHead( stage4 );
		clusterHeadQ.deq;
		let ch = clusterHeadQ.first;

		kmean.clusterHeadIn(ch);

		if ( stage4Cnt_2 + 1 == fromInteger(valueOf(PeWays)) ) begin
			stage4Cnt_2 <= 0;
			$write("\033[1;33mCycle %1d -> \033[1;33m[HwMain]: \033[0m: Relay 16 cluster head \033[1;32mdone!\n", cycleCount);
		end else begin
			stage4Cnt_2 <= stage4Cnt_2 + 1;
		end
	endrule
	//--------------------------------------------------------------------------------------------
	// Stage 5 (Data Receiver)
	//
	// This stage receives status data from K-mean App
	//--------------------------------------------------------------------------------------------
	rule dataReceiver( stage5 );
		let d <- kmean.dataOut;
		if ( d == 1 ) begin
			$write("\033[1;33mCycle %1d -> \033[1;33m[HwMain]: \033[0m: System \033[1;32m finish!\n", cycleCount);
			statusCheckerQ.enq(1);
		end
	endrule
	//-------------------------------------------------------------------------------------------------
	// Stage 6 (Status Check)
	//
	// This stage checks the status of the system and relays it to the host
	//-------------------------------------------------------------------------------------------------
	rule getStatus;
		pcieReadReqQ.deq;
		let r = pcieReadReqQ.first;
		Bit#(4) a = truncate(r.addr>>2);
		if ( a == 0 ) begin
			if ( statusCheckerQ.notEmpty ) begin
				pcieRespQ.enq(tuple2(r, statusCheckerQ.first));
				statusCheckerQ.deq;
			end else begin
				pcieRespQ.enq(tuple2(r, 32'hffffffff));
			end
		end else if ( a == 1 ) begin
			if ( cycleQ.notEmpty ) begin
				pcieRespQ.enq(tuple2(r, cycleQ.first));
				cycleQ.deq;
			end else begin
				pcieRespQ.enq(tuple2(r, 32'hffffffff));
			end
		end
	endrule
endmodule
